pll_m_data_clk_inst : pll_m_data_clk PORT MAP (
		areset	 => areset_sig,
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
